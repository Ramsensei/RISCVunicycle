class RandomVals;
    rand bit [0:63] val1, val2, val3;
    function new();
        
    endfunction //new()
endclass //RandomVals;
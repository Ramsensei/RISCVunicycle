module ImmGen (OpCode, InstructionP1, InstructionP2, Imm)
    


endmodule